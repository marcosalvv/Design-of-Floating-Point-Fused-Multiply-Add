library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
-- VHDL 2008 ONLY

-- A leading one detector circuit, it determines the position of the most significant one
-- Version compatible for the single precision FMA
entity lod32 is
    -- Not generalized
        -- IN_BITS : natural := 74;
        -- OUT_BITS : natural := 7;
    Port(
        in_lod: in std_logic_vector(73 downto 0);
        out_lod: out std_logic_vector(6 downto 0));
end lod32;

architecture Behavioral of lod32 is    
begin
    with in_lod select?                                                                         
        out_lod <=  "1001001" when "00000000000000000000000000000000000000000000000000000000000000000000000001",  -- index 73
                    "1001000" when "0000000000000000000000000000000000000000000000000000000000000000000000001-",  -- index 72
                    "1000111" when "000000000000000000000000000000000000000000000000000000000000000000000001--",  -- index 71
                    "1000110" when "00000000000000000000000000000000000000000000000000000000000000000000001---",  -- index 70
                    "1000101" when "0000000000000000000000000000000000000000000000000000000000000000000001----",  -- index 69
                    "1000100" when "000000000000000000000000000000000000000000000000000000000000000000001-----",  -- index 68
                    "1000011" when "00000000000000000000000000000000000000000000000000000000000000000001------",  -- index 67
                    "1000010" when "0000000000000000000000000000000000000000000000000000000000000000001-------",  -- index 66
                    "1000001" when "000000000000000000000000000000000000000000000000000000000000000001--------",  -- index 65
                    "1000000" when "00000000000000000000000000000000000000000000000000000000000000001---------",  -- index 64
                    "0111111" when "0000000000000000000000000000000000000000000000000000000000000001----------",  -- index 63
                    "0111110" when "000000000000000000000000000000000000000000000000000000000000001-----------",  -- index 62
                    "0111101" when "00000000000000000000000000000000000000000000000000000000000001------------",  -- index 61
                    "0111100" when "0000000000000000000000000000000000000000000000000000000000001-------------",  -- index 60
                    "0111011" when "000000000000000000000000000000000000000000000000000000000001--------------",  -- index 59
                    "0111010" when "00000000000000000000000000000000000000000000000000000000001---------------",  -- index 58
                    "0111001" when "0000000000000000000000000000000000000000000000000000000001----------------",  -- index 57
                    "0111000" when "000000000000000000000000000000000000000000000000000000001-----------------",  -- index 56
                    "0110111" when "00000000000000000000000000000000000000000000000000000001------------------",  -- index 55
                    "0110110" when "0000000000000000000000000000000000000000000000000000001-------------------",  -- index 54
                    "0110101" when "000000000000000000000000000000000000000000000000000001--------------------",  -- index 53
                    "0110100" when "00000000000000000000000000000000000000000000000000001---------------------",  -- index 52
                    "0110011" when "0000000000000000000000000000000000000000000000000001----------------------",  -- index 51
                    "0110010" when "000000000000000000000000000000000000000000000000001-----------------------",  -- index 50
                    "0110001" when "00000000000000000000000000000000000000000000000001------------------------",  -- index 49
                    "0110000" when "0000000000000000000000000000000000000000000000001-------------------------",  -- index 48
                    "0101111" when "000000000000000000000000000000000000000000000001--------------------------",  -- index 47
                    "0101110" when "00000000000000000000000000000000000000000000001---------------------------",  -- index 46
                    "0101101" when "0000000000000000000000000000000000000000000001----------------------------",  -- index 45
                    "0101100" when "000000000000000000000000000000000000000000001-----------------------------",  -- index 44
                    "0101011" when "00000000000000000000000000000000000000000001------------------------------",  -- index 43
                    "0101010" when "0000000000000000000000000000000000000000001-------------------------------",  -- index 42
                    "0101001" when "000000000000000000000000000000000000000001--------------------------------",  -- index 41
                    "0101000" when "00000000000000000000000000000000000000001---------------------------------",  -- index 40
                    "0100111" when "0000000000000000000000000000000000000001----------------------------------",  -- index 39
                    "0100110" when "000000000000000000000000000000000000001-----------------------------------",  -- index 38
                    "0100101" when "00000000000000000000000000000000000001------------------------------------",  -- index 37
                    "0100100" when "0000000000000000000000000000000000001-------------------------------------",  -- index 36
                    "0100011" when "000000000000000000000000000000000001--------------------------------------",  -- index 35
                    "0100010" when "00000000000000000000000000000000001---------------------------------------",  -- index 34
                    "0100001" when "0000000000000000000000000000000001----------------------------------------",  -- index 33
                    "0100000" when "000000000000000000000000000000001-----------------------------------------",  -- index 32
                    "0011111" when "00000000000000000000000000000001------------------------------------------",  -- index 31
                    "0011110" when "0000000000000000000000000000001-------------------------------------------",  -- index 30
                    "0011101" when "000000000000000000000000000001--------------------------------------------",  -- index 29
                    "0011100" when "00000000000000000000000000001---------------------------------------------",  -- index 28
                    "0011011" when "0000000000000000000000000001----------------------------------------------",  -- index 27
                    "0011010" when "000000000000000000000000001-----------------------------------------------",  -- index 26
                    "0011001" when "00000000000000000000000001------------------------------------------------",  -- index 25
                    "0011000" when "0000000000000000000000001-------------------------------------------------",  -- index 24
                    "0010111" when "000000000000000000000001--------------------------------------------------",  -- index 23
                    "0010110" when "00000000000000000000001---------------------------------------------------",  -- index 22
                    "0010101" when "0000000000000000000001----------------------------------------------------",  -- index 21
                    "0010100" when "000000000000000000001-----------------------------------------------------",  -- index 20
                    "0010011" when "00000000000000000001------------------------------------------------------",  -- index 19
                    "0010010" when "0000000000000000001-------------------------------------------------------",  -- index 18
                    "0010001" when "000000000000000001--------------------------------------------------------",  -- index 17
                    "0010000" when "00000000000000001---------------------------------------------------------",  -- index 16
                    "0001111" when "0000000000000001----------------------------------------------------------",  -- index 15
                    "0001110" when "000000000000001-----------------------------------------------------------",  -- index 14
                    "0001101" when "00000000000001------------------------------------------------------------",  -- index 13
                    "0001100" when "0000000000001-------------------------------------------------------------",  -- index 12
                    "0001011" when "000000000001--------------------------------------------------------------",  -- index 11
                    "0001010" when "00000000001---------------------------------------------------------------",  -- index 10
                    "0001001" when "0000000001----------------------------------------------------------------",  -- index 9
                    "0001000" when "000000001-----------------------------------------------------------------",  -- index 8
                    "0000111" when "00000001------------------------------------------------------------------",  -- index 7
                    "0000110" when "0000001-------------------------------------------------------------------",  -- index 6
                    "0000101" when "000001--------------------------------------------------------------------",  -- index 5
                    "0000100" when "00001---------------------------------------------------------------------",  -- index 4
                    "0000011" when "0001----------------------------------------------------------------------",  -- index 3
                    "0000010" when "001-----------------------------------------------------------------------",  -- index 2
                    "0000001" when "01------------------------------------------------------------------------",  -- index 1
                    "0000000" when others;                                                                        -- index 0
end Behavioral;