library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
-- VHDL 2008 ONLY

-- A leading one detector circuit, it determines the position of the most significant one
-- Version compatible for the half precision FMA
entity lod16 is
    -- Not generalized
        -- IN_BITS : natural := 35;
        -- OUT_BITS: natural := 6;
    Port(
        in_lod: in std_logic_vector(34 downto 0);
        out_lod: out std_logic_vector(5 downto 0));
end lod16;

architecture Behavioral of lod16 is    
begin
    with in_lod select?                                         
        out_lod <="100010" when "00000000000000000000000000000000001",  -- index 0
                  "100001" when "0000000000000000000000000000000001-",  -- index 1
                  "100000" when "000000000000000000000000000000001--",  -- index 2
                  "011111" when "00000000000000000000000000000001---",  -- index 3
                  "011110" when "0000000000000000000000000000001----",  -- index 4
                  "011101" when "000000000000000000000000000001-----",  -- index 5
                  "011100" when "00000000000000000000000000001------",  -- index 6
                  "011011" when "0000000000000000000000000001-------",  -- index 7
                  "011010" when "000000000000000000000000001--------",  -- index 8
                  "011001" when "00000000000000000000000001---------",  -- index 9
                  "011000" when "0000000000000000000000001----------",  -- index 10
                  "010111" when "000000000000000000000001-----------",  -- index 11
                  "010110" when "00000000000000000000001------------",  -- index 12
                  "010101" when "0000000000000000000001-------------",  -- index 13
                  "010100" when "000000000000000000001--------------",  -- index 14
                  "010011" when "00000000000000000001---------------",  -- index 15
                  "010010" when "0000000000000000001----------------",  -- index 16
                  "010001" when "000000000000000001-----------------",  -- index 16
                  "010000" when "00000000000000001------------------",  -- index 16
                  "001111" when "0000000000000001-------------------",  -- index 16
                  "001110" when "000000000000001--------------------",  -- index 16
                  "001101" when "00000000000001---------------------",  -- index 16
                  "001100" when "0000000000001----------------------",  -- index 16
                  "001011" when "000000000001-----------------------",  -- index 16
                  "001010" when "00000000001------------------------",  -- index 16
                  "001001" when "0000000001-------------------------",  -- index 16
                  "001000" when "000000001--------------------------",  -- index 16
                  "000111" when "00000001---------------------------",  -- index 16
                  "000110" when "0000001----------------------------",  -- index 16
                  "000101" when "000001-----------------------------",  -- index 16
                  "000100" when "00001------------------------------",  -- index 16
                  "000011" when "0001-------------------------------",  -- index 16
                  "000010" when "001--------------------------------",  -- index 16
                  "000001" when "01---------------------------------",  -- index 16                  
                  "000000" when others;   
end Behavioral;